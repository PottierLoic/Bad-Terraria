module main
import gx

const (
	// Sizes
	screen_width = 800
	screen_height = 800
	cell_size = 20

	// Colors
	bg_color = gx.rgb(153, 255, 255)
	dirt_color = gx.rgb(102, 51, 0)
	grass_color = gx.rgb(153, 255, 153)
	

	// Terrain genration
)