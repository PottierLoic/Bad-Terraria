module main
import gx

const (
	// Sizes
	screen_width = 200
	screen_height = 200
	cell_size = 10

	player_width = 20
	player_height = 40

	// Colors
	bg_color = gx.rgb(153, 255, 255)
	player_color = gx.rgb(255, 0, 0)
	dirt_color = gx.rgb(102, 51, 0)
	grass_color = gx.rgb(153, 255, 153)
	
	// Generation
	world_width = 50
	world_height = 50
	chunk_size = 15

	chunk_full_size = chunk_size * cell_size

	// Player stats


	// Enemy stats

)