module main
import gx

const (
	// Sizes
	screen_width = 800
	screen_height = 800
	cell_size = 10

	player_width = 20
	player_height = 40

	// Colors
	bg_color = gx.rgb(153, 255, 255)
	player_color = gx.rgb(255, 0, 0)
	dirt_color = gx.rgb(102, 51, 0)
	grass_color = gx.rgb(153, 255, 153)
	
	// Generation
	world_width = 10
	world_height = 10
	chunk_size = 10

	// Player stats


	// Enemy stats

)