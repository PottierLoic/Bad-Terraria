module main
import gx

const (
	// Sizes
	screen_width = 800
	screen_height = 800
	cell_size = 20

	player_height = 40
	player_width = 20

	// Colors
	bg_color = gx.rgb(153, 255, 255)
	dirt_color = gx.rgb(102, 51, 0)
	grass_color = gx.rgb(153, 255, 153)
	
	// Terrain generation


	// Player stats


	// Enemy stats

)